ENTITY DECODER IS 
	PORT (        
		D3, D2, D1, D0: IN BIT;
		SA, SB, SC, SD, SE, SF, SG: OUT BIT
	);
END ENTITY;

ARCHITECTURE RTL OF DECODER IS
BEGIN

	SA <= (((NOT D2) AND (NOT D0)) OR D3 OR (D2 AND D0) OR D1);
	SB <= ((NOT D2) OR ((NOT D1) AND (NOT D0)) OR (D1 AND D0));
	SC <= (D2 OR (NOT D1) OR D0);
	SD <= (((NOT D2) AND (NOT D0)) OR D3 OR (D2 AND (NOT D1) AND D0) OR ((NOT D2) AND D1) OR (D1 AND (NOT D0)));
	SE <= (((NOT D2) AND (NOT D0)) OR (D1 AND (NOT D0)));
	SF <= (((NOT D1) AND (NOT D0)) OR D3 OR (D2 AND (NOT D1)) OR (D2 AND (NOT D0)));
	SG <= ((D2 AND (NOT D1)) OR ((NOT D2) AND D1) OR D3 OR (D1 AND (NOT D0)));

END ARCHITECTURE;